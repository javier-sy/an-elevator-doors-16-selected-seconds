BZh91AY&SY��.DqN_�ryw������?���  `��B��D�R���� T�BU���P   (         �  h        X ���D�G�:u�Zn�2��ݝV���ܻg'G�:����w �ѣJ�:h�Υ��FCA���G ���uN�D�E�ZqWv4��3CMr݇ k��@����9I���t��t4�M��  N�MP�ӫ��`a�N�i� I�,�.í tWAݝ���N�����S�v3�� (��m����8n   d�@���h����t uM`ínç8(1�m����5���ˁ���۠a��   ���:�XCFF�M`í:gJ()�v
t4h�ʺU���CGA�:|QD�@"��U%P�~`�J� h  2h�h   ��!�J�(h0��0 �0#A�"��
��2h����0 &�`���eT�
���C2 Ѧ��a2`�$hL�L�M�<�ɲQ�4z��!�=&�z@I�Q
22MMO$~�➧��6��P��F����ʗ}��=�Lr�w�I$�g���BI!��BY i!	$�x$�Hc!��?Y����B�Htd����%���������;W��m�x�{�ݩ��w��5�:~���wC��@!Nف�`�(C���,� BI �O5�X]��S�ā	$��C��=� rm�y��F��zqŇ��2�y�w����C�#}L)�^ϑ�lYg�/G�+�R��{�e!	$���kɯM�o�{)��oC�(��H���ɞ|rZ������}��zs��n�9�6����-�
�����n���LZ,{�70�
/b��o�Q��`|�X�����.��ˋ[sEܩ�<�qe�WA�3	��d�V�ƪ$�ѱ+f��f�u*Γ�qOv�+sZWR���D�����%ђ���0Jx����;EI0�eVff�H��������K^,�H�6'�[�Y�m̽3-0wbS4GX�PdaQ��u*�	��*�b�d�z�&mc�p��:��n�E=QFf�4LI�z�qZ!��̶$�iĉm�f5HkQa���>�J7�jJa���1h�0�w" �+&���{�����|��wJ����9��wb�m�7{[V\��3V�Nڻ�6Z��ɻ��Bi����1LyB(k�1�u�Lȋۡ��B%Ī�Q�Ĳ���؂`_����O;CwB����f��V���J�1���l2-�hD�����wKK�~0�F��,Q[U(�/.ԕ6Y�4�B�[d�ea���Si�s-Q���Yy�rSCj�D�Շ��Ò�,��!u/�o6�M [�ROT�Z �8���e�w�."o���1�Y� [�
��xk귒\�(tR�ɸoT9�k"Օ�F@��V�ؐV�
��cP@l�*�;�)S�X/t,2`*S
���S(���kǂ@����]�ܭ��m�2Lca�.Q�
:�k�P.�3��A4�X��%��6>��&�k�D�I,d����3-���{@��j���Ub��`v�39����D�ږ�D0�����#��iE�'eb� �4��Ѝd8� {�#4�	��q�C�R�U��^��¤��ՋE#�h�ݒ�:(�Ec��i� ~�S5�9 �]�& �i��s3b�X��&ɚ��{V����|��ˤ��%�����w��۲�����H�d*�T6i��q�|>�`�b[9��h�εq�c$��wr�A��R�V�b��G)���s1XÒ� +v�&�j�ř/T#6��f��ۄAw����6��5�Www���)
c���G�1�^Z��a,FP�{���Ֆ���b����l�Ȝ8��ld/ay�+��7�q�K��F�W2GAk������n��3n�[�(��f8h��g�^�x�9�^/�n�WO�PP՗F��$C�J�6��%�x�O�pL�1��w[(=���f[��@�T��;s.�͹��뻡�EW��[v���Ԭ�"��m+����*��˒��0��'v�"��މY����Ѻm0+��w"-��ʘ�X�%�iV.�:u�1*]S�5��Wv�T�HS�K����X@�n�(4���:�a5h�z�lJS�ASv�ˆ�Yp�A�0dbM�e%����m�r-��`̖hf��=d^V�$V����F�˺�
[W�C ̎���n񛭍MRCfT���\�Y����fe���q`�h�2�ue���M��J��j�zcPB�ӃH�[��#�L�-m���ыi*
��&[�S1��j�B�/�J5d�^��v45m��7S�l`X�Z�;R�A�L��)�d��b����zo.�M�N7E��=um�͔�E�Ů��+X�?�Y� ����c�kk(��-�*�j�Z{НSn*�f���k`��5�)���^�w� O�-� y]^�KcW�fi�$9t+R�R����xM����6�jS��ڗ���i�p�i��q̠�I�� �p��+��k��o.�h�*Q3Jb��2Hu3�e˴�m����Z�3#��F^B��Tڲ�0�uJ%Y�{`�)�Z� ��"��v��)�@+R��_K5�-S5���0�ԭ�z���a��MC���4�[En���iYUSf:ɄZ�j�nS̩��6K*�2�e�b�nc4��ƍe�ֱw�z��<1O�"E3�3d�%��t�ln���m�h�R+&��F�U��:�Mh�YKi����Z�e��W��m,'C4n�Ȅ��#-z1ә��5�Vڸ�y�R��R�s/^�]RjP�ƊZ]���m,4�V�O*� ?e�eD�"��e*HbN�֗4D��D��)`H�n��鬡y�h����ՓZ�ݶ�j�˖�|�Yڴ,CYeo�5��QAc��m4X")���~��v�2cy#�;p� �,�F�cT[ּ �U�^:i���]��ݕ�kRy�̋0ޤP&k����f�;s�)	 ��uM{t�Yb�`��j/���k�%u�6��u���b��XΈf�M�n�ee�.S�Eu��D[g�Z*z��KBkU���&�~��-�Vk$\�R�4q�fH����]�h�f���d�i�Jɑ*� �2��I�uv ���C���w˭��ƌ/jm��ֺ�))�ɡ.^d7x찦�N*sXst���B��^�w-i��T�,��ec��Y_�ff5�*`�[�3H�f��ҥ�{P��cy�K j�y?iW#kT04�i{�m��Oa��aM�ܙ��j��,yY0�5�n�ZZ�nⴆ�7+^�.���lց�);�I@;�kJ�+>���w1��W���X�u�0(���(��=��7KA�X�fK+A�Q1N��NJ�n3��.7����Xj�@'F�x�h]�5��;yd�j`o3�V�R��
S�ȭ՛Q�+l�׀	��jڦ+f�bTvl��+���>�U?��}-���ֵ&���M��љޜ{ۻ=�d�awO����]��Ξ��ܼf";�\��]o�a�:EsZ�09ls��W�N�ƃ��݉{�����W�g��=�Xn��v+I�{�d�,x�x�M��.콨��.j9m�J�j�]V�FѺ��)���ȒB���d��z���^:w�=�3�n�n����:6�=�:I����,Y����rQٻn�u���>���::;��tv�u�ΰ������\�qL�u�k�����hp��Z,��7)���QC��A�5���l7n��;�m<	\WN�{=-Ӷ�;t9��]��s�8��/�[�ۃ��u�hC{�U�&3g�d�Ѡܥ㧠�d�g6��f��]�1:%���Iz"��];��q�;j�Ѻ*�mk�ohWX�#p`|�N�D���tt �1�ۺ��l]�<ٹ�-�Í�up��	҆��qlpM��ćm�w�ncn�8\֝��lu��.��r\)�S�^�o[�]����?1������O5�8��rY#ܶj9Խq��x��;�q����1I΃tn��'\��e�1��ԏ��,�l�i��8^��հ�]%H)���ٞ���\sk��*�2/Fne����]��j'�q�ۍ�ϟ:E��.qnb�dFf�SWq��3c�9���^y-.�I�u�۳����tQ����95ț������^}��v�w�Z��/n7.9�c�";q�A�}':�ݺL$:�Y�H��Qt>�މ���7iZO���L$�k9�3/;q��.��\��ݎ�t��n�����M��= ��v9����䱼�s�
��\up۳b"K��Ϋ���t�݂�]�G��6��'V�V7�����/\۔��v
��n�F�����u��<3ݽn��q���7.� �@v�n-��R��l'D�\�n.���`ŒԹk���qζ���g�裞˞ìX�/���b�S��n�������]�z�8w��w���$�[�M�Kt����jm��u����v���;�Z��[sٍ�6�琼Ƹ�M�F����+��q�'5@rW��aI�9ׯ{F�n�8�Ld%�ݎ��=m86��Ǜ�n;{ǔ�G��c�ٵ'Y:NM�����͗j���Quv���GT]�y�F�펳ÝJ��r�]�� �v�Nn�ٴ�*����m���x	嚷���ݻ�oG�aΫkS�k=�r=�9#�ݶ�^�챻j��x�h;��^;Is�ٹ-�m���[uX�z�q��F��m�㲝��끷n�#�X�2��M�[�.�ǘ۰�6�*u���`��s��e&���Gsv�:*�/`&v�v0���Ź�� ���~S,�۞=n^�cGf^�$ݗq�z*[���$����\�q��}d|��S�Qn��[mQf5�9��k5..�+�1m��'��æ�6�$�ܽPݝ��]q��tn�s����v�>!y;�]�u��8�X��m��&6:F=%���w>:�ƌ粰�Z�ql��O���ך������vz�X�r;�:z�U�;p���|_�e��m-��v���g�v��8���7��/.m��'s�\y��	7mK����H��LgnM�[8�ű���r�b^�t���x��8��\�v�/�iv諔R�g��N��X�vՍ��u؋����tO��nL`���R٤S)�]�AV]�]�hٹ���]j�r��;p>r�yC/n�u�utn�]x�+���n���۷#e�T�m�=�����P�v�� O�c���7q�Y���5z�Q�������n۱���m��q��ku�G��6tl��F�E۶�7��p�4�ݜ�Z��㑐'��JغF��.1�L������nx�M���+6�4���:�q�m�Vc�(]�1��p�؂������u�8P.�k�d��]�]V1U�/e�kO���EY�71�n�ͺ�m���������G�I!Ǯ_͐$ 	��e�ol���Z:Ng���w��9�iGճ�����������u��z�l�(c���q�x,5��<sMV)8jT�++�ߋ:iYP����Q^�.�F�3
W�|�qצb-gl�F���ì���8-
�Z\�2�a�0���,i��J�m:8eY�4����km*�)�Y�V�R�R�]ut��R��e��^Zb&�m�
��a1y�'km�YY�WR�*�M�eL�¸�TEQU昊b��ÚQeTkA�K�J���k/q�PK[c*���ZmmQ��J��iV�뗇C
ѭbSEq���0̝�)��&�p�cm��Dn\N�\���5�ņ�[I��eAQDm�5�J	j�\��	�aE^Sr[J,w3PsxÄ8���d2�3J��H�Z
�TiTT���g����6�Ïae�|�c��Ps&L�fcR��0���f)�0CV6�UC+J8��kj6�iҜ���U���o.2�ek��Ѻjbe,[l᮶m�m�J
���f0�l\Ze̖�ƫ�2^�;
��mF��7q-��Z�m]��V�mbms0.\��*ԡYD*\ܩ�׭3(��[EZ0m�VW�J�ۨ��T`�2�^���j�m�2䠮��*�2�YAv��R���1�*0�ت��hM���a�V
�,D�**�᮱U]u��h��D�+Wܥ�)ir�& �TQ�Q�Y�SZ�Z5�J��Q��(b1��UH�ܪ&5�l�[faUb[UTX��F#�A��r�j�����*���ҡX��Eb�YR�@��KHڱJ�̰+�YYX��!��v�:�,U��DVÄ*�8h��LIX��,�ƴ�**�V[B�UT`��-+!�Sd*��<[8xI���Ì,�"��+԰;$�q���Pĥ���
����AA`��b�-�Du�ڋ���B�aY��0QIm���,\eH�+PX�aXLf$Y�b��`�e��E���&�

�X,UPX,5
�j
ʄ�Tm�"quYH*�q�[�H�H�� S�0d1�������%���(��`�ac T�)m�d��b��E���1��n4��`����
H��,X,UUee�`���Ȧ��U��
F"����c*�`���E ���*��+ ��UE�H���XV*��̪�`��o9�ANx�*Ud�ذR��Y�������,kCTR)IP��R�B�eAE��V����/V�Q��F�EC���*)�`�%dDAX
b���Y�r��B,U,�,�ҵ�
6�1��V,X�+%�"�(�c
�b�,�`�F�Rm5���$D(EQLjR�Z��B����E��kYY-l+���]J��!Q���B��[*(�cU��֎Y���k-
�2�X�T�5*E�̳�V�p��
�V�T�-+���Z�Q��iŒ�#�^hp�Rj
��L���u�J�-
���Km�[�LNm�¥#�Yeeb�!]`Ua����j�3r���rآ

(�\a�R�D�+�LeԺ�q+���e�hDFbjL��	X,���w$111+"�n�V�)����HbV�a�r+�!�H((��s�LM���]d.��.a���-��V���� BI ��%+����ߏj|zV��pE���Rp�p�q&g��_f4�����v�WLP�G���sf���c�r��*z�����8��݅��L����Y;V�od)�6�O6^P�r�q���kg��'/R��2�q���nS��ۧ��s�:@�����p��|��]�r���{v��:����{[�rY�m�ۭD˙�i��˴��[H�C��qjݘ-���c$u�;N1.������k:��;Y�^\>\���.�[nZ�*��i�ۓ��C��ƚ��G��M�ln6�����:m�7m���Jx/n��F݄�����:U�J)[�݉�/c'��<5)V��1�m����p��]sn(��z�tTh��hr]s��vOny쮺�z77���֍���.cs�3�"��on\D��]�z����d,��[��>w��܇w�����|����U�چ�u��]U�p���ݰ�<�݂3K��T�qM[��f�uZ�]�qx�'<9��K���ocK���9p�[�1����l���nf#m��c�>��<M<�s��݃�w�w�J�����oՑ�H���^���n� �X�S�,�y���3�b����uu#8p��.��+o�{@=.��)>��÷�M~O������[>�~�ꝧ�.I��lN/�w�1�Y����k����D���j	bbH��I���z��dm��Ў�F�<�/y����4�>a����;N�W,���w�m��$�Ĳi�E�Y��L�}ߤ�j ���-�K�\�Ξ\�F�cY�aT���OU�yc�U&Y�c(ԙD[�������C�};6�\�ݕڠWv��xfz<�)��k�|��	m�b��q�'d�"��A@�K��	|N]tr�2k���kx&N��I�C���H��79��4}ݵh���η��C<$��	�zK][�u�SYy� �����",�J�~[��ɇ'u��
�v�n��
o��Gg���P�э�������%Q9�\�/.�He�%0yX�A�Uu.�~|���|��s��Zu���d(n�7F�pֆ���7��]}.�X�b�x���,�	y�77�ʘ����v|&.�-�o���� ��+���Q�`Z�)�����y�!'f�6��*����~�s܏�>oǻl� [��OPT���4�h�ݾ�����o�����cv���i��`�-��1�A�ڕ��^����:N���FrK�6��j�%U��u%��]{�scL�©���}�Eih�݉�w-���*ʗf4_�f���"�."?lj���U+/i��Fs������x2��}w�u����� �� �����{�.�t}�%�MU���w��{ͺ3L
��Tg]s�HI��-�M�\�U��z3e�C�]gn�]�&F��t��a��|(��<�����q]u��w+��W�p�"*]yɇ���v�u��ug�������&�BB0!�
�2�l���5r	�p� �S�y�c��vBi�&$F	�����\�W���%Tn��	L0�����2�S��=R��z�{(E����KǦ����D�=��ײ�
���H��A�sq��V�SZM5���Mł�m�u=v�ӻ[l���k�^��=�q�+��:�;N�7ΐ���XF����+9�	��Ҏ�9=�+��#W����M�r8��64���!����4�U�T��9���,dU%eD�N8��m'D����ѡ{�z�ǫ��4��	a��<s�~�w����u��bu[�[Tv�kq�٧x=�"4�us����D�z��>o����n�6�����E�@Y^6h8�j'�7�P=��hc��/}��y�(�Eo:��s; ����i�޿���5[�L�t��8��_䷝
��
�ԺV٤x'i�Lt��u��1U
�h�7���Κ�wc�k�Ҝ�����������ߟo���9�nm�f;vܴ�Æ�l�ᅿ
W~����-Wν�g�KR���L^��!z�f���5�N��ؽ!\�%�Eѡ.�_VK�9��,t�VX�0YG��=�[�OL��n[�6�Z��pʵ����y]��P�v
tm��4�
rH�<cI��A�V�ʆ�lee���r*s5/���]�j���6�8Fh� XE��4�ɘ���L�6��^�om�E'��s�Gu�Q;��t�����~:�4،H��u{m�`{wnF�E/ce�;I��2�{E
�9���C�o},%N/{����o>���G�^���s/��1,�Gæ�������&������{Y<�G���N����\���۝��;V�<��k�qm���A�m�R���t��S�g��vmخ�S���pf�v��un׫s��f����Ȁ��_\]�i�7̎��䗍η=)9���{�������o��w��� �:�\�^�h�8��Q�:���μt��x�vW�8��u��k�]�{ja�@�����n&FFEL��7i�̇���}yc&��~�E\�*�^����#y�=�i^qGg���u�NF�����<�#l�c۾Q(j��L _�`�_�ݏ����"R\f��Ǘ��f�����jWnŷ�j�rX�oq�_��5�'����r5��M��*�
X2�ٲ2���<��z��7���G�-;�����{K��d������!��%b��P=#�?���%�����������u����.�.�WTn����h���t)s�E���g_E�����K��MLr�%`�������a���wj�}�o&ފ�ζ��㍓
���V�gu��=)vr�l��2�����j�j���fzP�������LD�A�x��nHmt�Zҫ��+�����9�T���e���z�-Ƥ+Q�*�t���N�kLu�Xi�]tTs�c���Y[��jc�z9�Jk�GZ�K��n�-6+��ŚEu�ȍ��j	�8f;� ��lw˛�L̑��9���4seo;6���l��Wu"[,S��j�ө2@C��8Q��=:�KdG������ƶ]v,כQ�ǅb7l&_Iz-r��r��*�Ա��6��u#�+�ƴ��4�� �/5J�$ӹ���^���~����q>��0��`����@�����L�E��������(���/���
%�[9�����?��i!�B�k-惂��L ���j�m���e�@W$K���!ku�����o���ժ�-�p�����}A��������A2�1�58'�bQ�Kzxݵ��[5���re/V��_eb�n�I���s�d�;'�M�eßu4�eQ���;�t�0=����h°8�U���n���hY]3�l[��Kj�+J��נk���u/�'}b�̊�ock��w�3����t���8~���n:&�����$�Ha�P#�D/F
���	���u��p� �k�N��6��B��N1T��Xt��ٞ�9� tv&:9����3@
� ��*a.^Lr	�F��c�� ��}�y���O�Vl��z���Ɍ[�	�(�9h>
W L���.���U����Q&��+�v� l3�l^d�� ���s;l�|���Q4]�4�)v%��'o�����`_-tvw0�Ŭu�]�n���
�gq˝��:�x���ܶ8�d��޲��ҹ8Q,�9|��\�>�B�.��<=�x��Pك����������W/�H�l8�a�ڎ��:�0Z�Dlk�?��3�W�ʧIQ�Ο�%��G݇2��gL���	����	'�r�7 ����rM$$3b�:�s[3��:Ux�5k[e�4�ݚ�PM}=;z1u�y�ό�ζ�A(7��L,��W���=�k�y����P1�*�_U�h<���f�p �1�����Y��`��˧Yy��ZڮU.���~Lf�jO��G~�*����Az�g�lN��+̪�.1�e�b�ş �C�����b�`�I��������ڎ+ܞ��^�i�A�e�~𡙫����z������>�� b�9�hg�tĴ",`��A�5�؜��(ޭ�y�k���g��ż���׊�I�:�P1�/o>(8D�ۂ� �1��B]Z�ݿ?>����~�����u"���崾�R�$*�V��K���1�Z��j��B���D1��X]�|�6�c�{eQ66	\{ݓ��WNu��4<�p��o��J��SHƝ���K>�u��P�F����۠��#s|����m�������m�T�6�����f�
����O]�e��}&�Җ��*M'�� �.��������^���{G̓O3×\��j�
%�I����'���U2��92~�l{p�vT�a��K�����U�}"iP���ܴdq&_I��uD}�70G����H��S�y���I�=XW��c"(������}�O{3��-'鐋�<�w��`����OayN.���4}��<�ڃ�++;{�,��w��7
=��!���w��֫8D�@��|����bA���	�.A�`C��Ǫ�͙��ﯣ�v�~~�X�ϟ�ICo�N��q�<���N�=�*g�R�b8�j��Ƅ�:�S_�T{!��g�F�y��V��wr�3��^��S\��T�~��I���Z*2��N�(UkK`��f'9�|�#�zym��pM�i�UVF���,̶����Y%�8a�S�<�;��XϽ����6�P��l��9E{��ݥd�P��'DY*ιy�v�����<$AZq�������C�n�b�nY���G;���9۔���z�n�Z�$��ۮy7E���k���'a�貹�"��V7������e�ӷ�$"@ބh+�g2�z��O������+��>9��ǳ�%J��R�̷�Ȋ��R=��p����1_�C��'����uP����?Q��^w��6�?|�	�r�6��������)B�.��ʖ�f�OQ��`�H�7g�7{Lֺ���U�H���f�}�Q��Љ�����z{kS��:��\�͟���bsT����ȡ<b�=���a{T�Pg�/4��%Mbw��������k��m>��7x�j��y�xP�m���X�3ʅ����e�����̝�?P�`E�������8��z�ӓ��k�H�����*o$��F�mǰTJ hK<�y է�×yyS6��(C�>���}�[��K���� 6��{��Y9OQ�~o�߳{9�3�;u�v����l2R�(��Ι��8�{]х�*Q��F�U���$`�C��[�^�:���_U?>7&��пԾ�r�$�;�A�5#��Ĥ��0�%l���
�0"����:�IãI�XC�͎F(m��T& �T2�c[� �Q��yf�"ycg5Ez0gr���Fn�V&1���V	���d8�<�N��0A/�YJ%>���V�z��>�?�w�͎��M���#`Ǎ��,���Ӕwdlk�z��a\���w���k��q��䀩U�y0��뺰��WiϢ�8�Mą��6N���"7���g��Ii���K-fZ�7�����!�?=7����c��ܾ�+��1.�m�e�j�'����o?2����v��=�(`�>�z��[�y>�.��|*O,$�?��ۚZ�uqs�]�E�5�J�D�η��4G�����"hwr�0�`8��x
n7��g]}u�>6 ���hr'=׷>�i� J�dNg8�����������o�\	���@(���N�
7�
c��ܟ�[ɡ��X6b�A~���,� [@M3B'et����9�~�Q�P��}��G����"'�q��1ug���J�b���r_��F�銚5{y&N"�`�M�L��p��Tgj���|�T�ۮ{��a�����˲�����4q엸�tR�����ܪ��כ�#��:i�<��R׭��D��j�b�N�Gj´���)����A��ı���᭔e]�.�WR��#xt�[|B�^��X��w��ݩeN��Տp$����s�|�v��%�1f�9�h���Y6���B&��r����6�r�ͥN��oY&��U�=NX���ZS�J�G��V��a�+��Ks���Ν�Uu\�W���N���)���O\��\;��kZ�'mctF�˻qڬ���XU�nz��n��ۄ=sÔ��<a��k�W;p������X:y9Ywg���X\=,8�y؃��;/C�=c���l�i{u]����	��G���w{mԡ�����+gv����۠$��x��0�ң��\Ou��q�_/�$;p쉉��9�ۣ����:���0���ӤMm�msc�N{�ۨ��Ǯ�F���ֶ8�1[�k�7�m�jk�e����T�\�p�6�O.��ϑ?<��c�B�c����G\�n���n(�[\��Q������s�q�J���{��q�i�Gn�V�eg��-�DY��P�.�.3�=�yj�Y���qp<v���bH��3sZ\�Gr��>��(Hq�Kӡ�=uŕ3����!���.���CqwFP�Ukm�K�S���:��<w\�pɍ�m��\쩊���絷�vGgq�����6���}5��|�W��O�*�/����ߕ��_l��]���R��ܖ���mm��ˮ��u��+���I4{Dp?��m��9�߇�W">s�~� �2�E�Rk;jAkI�䩠���ڕ�1��xn,\J���'k����
���"D�)΃�gU�x����,�"pf�o�@��\����# �C��l��ۋ��_!��*�l�x��q�ڦ.[���������]@_P(NY�Omx��/U�oV�����Pk�v��P�Ѿ�ԉ�3�N�}�ߊ�+�G2�<�kG�|K(A^���o��(U�vZ�aB�8�tX�k�
1����6������v�����kw� ��71���`
�s�Ң�.�z&9�F}Yv*��(n9MY[���}�|�1A͕�!���~�ϯ�߷����cv��F�m=dZb	6�eTH����qez�i���2v~�h{�����B��S��|�<^��[:� :%MG�o�V�:�Xn�������c���t�_r�M��탔]�T�c� �5�M��������طm(�����G'vFF��@h{ˋ���y�u|�efc�u�c�m�d�q�2v܍������,g�8�j�t,7�9���Ѩ�_
��F"�K�44��s�ߣ�����!M[���2�{E`�� }��ĔWj�HI^@u���;;���ƃ��9�C|�y}�}�1�*:��H.���r��%x��yY�{_���~Rְ��n�kR+TA~,V���m?_��6����0����:��?[Dҷǵ�ѦQ �fK�H[�Z��B�!`{��G�G�^��}��J�V�t�%�J|Q�
(7����{�3��Ĺ��(q���砪f������v�i'6�M����]����O7C�^z�IX��Έ���g7)�v��V>�!��|��]�+��+�ǷA�$D+'�0��U坺�=Lq�9��=[��h]J��K�~�Go(���ڇ��Q9SÕ�9&��*��.���� �q�^�ჽ��Ɲ�;�CiR���W��]��8��Q�y3���������w���k���� }{&^�Z���C�f����E�����gj��]�앶��<��[�s��W&�N�Ms��׎ͭ�����r���g8��Hq�u�]PIʫV�֒����rn.
�&�_��+M����^�4�o 3�� J]��qq�Pq��_[5�
'��'ל��8���@����>�\�7��<��W�T	Y�,B?f���G��ެ��<�N��I��̝}Z��+/i�&�g�D��y.��Aݪ\YRN��Ů˧B���@�7�X:�"�u��u��Z�i��AV���ɫ�����N
�QJܲz/�˔
`�y2�o�b��Њ�[g���]�nT۾���'�T�=E�BV��{�,U�zH(�[�&f�s��N��R��$։�z+%F�4����Y��=�ǀ�V;�s������Їa4kΎS�_�Qz�������t��d�6 ��x��K���<���c�4�i���X��"����p;GC��i�3o�}���������R�,/T���__̘���.JY��s�U�'{�u��;��a痭�R��k5sήw�!ޡ��{Ж�Z=��0{nh��r߈!��Gp�-��R6��z��X��g������"��;\�B�>���
�h���hG[D����z�hCw3!����)p6�l�Rw�����
��Z��=�>�_����׿~��n�nW��H��7.ɇJ��,���OS]���LFm�0d�+�c��C��8-W�P�H���0�drH�5`�nVlfxu].��bbdȺ2'm,���VPdm��`�O�1�PŰ����@�Zj�ǚc�D�O/ ���ϫٯĬ�߭�O2\c��ޭ{�S�r��]�@����A1��Z�izGQ��9�*�T(�7���Z��������;�;Ђ���|`̞��O56��Q��^��8X[Ҹ�IR���~]�aD}�|����$o,����7��|"֊3b�w��Q/y�2Eфc�$��c��W$�����b|GBm@����ۊ������$�m�\'3ʈ�pݵ7�԰���F;I�󅶥wқ�=���y6jZ���,�|Ɏ웛!��h�p�sk��Y��|���TU�F{m��Z<s��غP��m$���I��n{�D�`�n�۶��ڻ���;��8�c���q��n,M���W;N�B�v���c�q]s�Gz���S��4���_���}�~}8,���ۭ�d��������d@f7V��˱ۥ�!��� �qx��C<����U*P�T�������CG
u9(@�G��ঊx7�*�z��Ɂ���/T�k�=[e{�607}�N�b�i�xQ�Gc�q!YZNq���TK�,�P��`6�n��8�d����~����w�-�����\���~~vF�Y{F.N���@��b+m_���}���w�ۙb�T��e����$��\��=�$TUaS+A\���8����kͯ�g�2a�C'*�^��"	���b��U��/i��zo�}�/В(ȩpGԬU��<	(f~2%v��%��=E�y�A��O{?L�|�K���6�;�%�ghX-�q�U��Z���\-�޾�R�+�}5�P�.�'�oA��b=�Èn�gi���.1.8��6v*��Xڍ*9��J���J jƫ�D>�JU����D�w"��g�*�T��0��Q2#]�� �i��7aU�L��#�VeX��e� 7�u�.���5R����ze���q\�}ڜ��ǻ�\��i ��|2IB���(u:pgN՝�:��{x�8v���Z�������=&���}���"��ԳG������.J��:�n�gS<���3h�owӗ���v]��C�-f�� b�����y�+o��qh�F���oޫځ+��0x3�4�.#v��]nOh���u��6
��������m%���F�!W�F%�/P�w�G�}3^���\�q�[@M��d7~ޖ'\%���2�?f��諥Ƚ��Bi%�s1�Ik6�-�%+�I|���M��a�6o~k�`7�q��[�\��,�ӷ}yt��h��Y ����֪�\y)A��5~��lʞ�>]t�GР��ɅִUA���5���y�L��Q �,�gK�J�?lw�^�*x�����ZH{`Z�+~"ji���-�w���C٣�����Ǟ�=�m%+@7�UM�S����z�@�Q'ˡ`��}�z!J�\�+��\+�~��~|����gpw�K.�:�GJ2�m&���,��	�}�o4(_.�uT��N�F�ypM�{�Kr
Gz.�Yo�ȶv
d��CP�{�C���gn�L����slP���1��>�s��9zՉ7��-h��tO��xl��O&�qAi.�=q'٭$��^>���fꉬ�����'�mPeB
�����.&%h2=A@\C~/�m�����{/��s����|�NU�KWm�ckK�;�cT��MӬ��_>?#�Ζ�r�t��Op��F`�KiEɣ/&�N�{4,���p%�q�b�VM�yz��Γ3�M��\_��8����?5}�?���D�}�g���P|��R�����
|r�T�&���0ǁf�S������E�Q�����M}�� �q-t$#1%�6\O�ϸs�d�,�'�1fj�/.�l7�qs��� M�΀�*|����W�ܑg�^O���5����Uk����!(PE��89KSj�����������)5��O�eYqY�n���jxڌ��A{�ǯ_	��뙙��E�Q�N(Mx�5��FOr$g����:��r+咕3��f&���d�I�}�o�����=��,���7�h������;P|��Q,�JA{���5:=��Ǆ��1��v�M�"�|��/����E�B��ß <�}#al�dJ�Q ��L������[�_ӱ���1Ï+Dq�q2�eU6U�;�&�.-+)�Ѻq���'I��c\�TV�z���eLT����je/{`��3b�����;8�^	���L���ڥ:�{�CS*2G,Rխ_9�]�R,*����*&|�gf�W|7�'\6=%��w���ݞ�����y�K,����6�19��X���1�SPP����߯۾������w����<Ť��m�����,��W�@������Y��_r�����$�0rY�.������`�)w��[����,md�݀ӥ�(��P�=�A�J�]
����<	�0�Y���ՠ�oӆ��v��i���$�w�.��X�����hCb���=Ԣ�][Bخ�;biؽR�@�'�z��	z�԰ ���؛�� O\g��9��v5�������ڑ{/c�\pyK�Y��L��=����z*5J���*�w���e 0�~5ނҤwB��q^*+'�I���|���"2{ �Zzp�~��2M�����꫍o)��T+N`ɥ��J�5��y�>K� ��̀}Mt�r};9���+J�G!9SQػ�����ib�5�P�|�
�o���P��>��Z�㇏	z��.��v���Hr�d��J�vՒ�(�I��q0a}��]�k�C[����]]��ή3�2��:zNG�M��&ᠻ4�n�!�va�'A��1"i�֡������������w��}�=�ZsBm("bs�4#��ڂ�6:��:��t�#��JO��l��fOh�:.3`\4����q��;��K�b����6G^(�I��Ci���nԦ����8>�6��,�1^Y��P6�f��k��~�v��o׺��{��JĠ�樜�wYE�K��q���k=^tv/����:i�c���E�S+H���Ý�]����F^|,��Y���<��j�{$8nB�-�$������4�`����n�8ulX&����0}�� ��zL �s1/��6|@�:��)O/�Q�`�o���ɚ����y;t3���3�V�|��&㘅���y5��ٹM�x��⠘�h�0�t�a���ѭ|�N�]��"�W[i�.�`�@VhD��&<OA�������F���@m��1�ټ�P�#�R�ף W��6�yvrty?;�TD�n�52��z�m�fų2H�Za�Y��T�����ۯ���eZ���g����V+�h�ny��S������8�XZfT�PL6�앓�Ec�oyzhF�&���1^؆'�R"kY��&�R|U�W1���}�0	�z���F��7�~}�ܟ�;�O������P(MAXϙ�:Éѻ�C`��tw���T$,��Z��O�d����UP{ckH����A���jS���z/���S����K�&�<i�j�`�J�~�N���I��P�=ܤ'>ؤ�N�fe�ۘ�nnViN'j}^��@��6x����I���d��{N��:�����]0h9k��#�}��D5���klU����	�B�όʙ�z�hf"�v+��BZB��52�>�#	8��~�G
:�$��Ƥ�؟1 �'іNl~�7]Q��%!�Ɯ�A`��3��x����*����$�.��#B�R+R5���ލǎǸ�f�te�x!��Iϯwg't�b��$~#�2b=�z��FtwǴ+b2�z%T��@�F�����܉L췆��KWe���x-B�R�5�sy:#��r��'��{�*������/"��~�sVB�5���J�:�E�T%��ԛ֏o^�Z�IO9#�1aR�v�C)Pε���I�fdx6�ҏv��:������&�2$�]l\1e�'F*��+kksWo ��jΠ{#;�F[���^`i_����8V��╛M�V
�|:<޻�8��M̉��V��Ǵ��'.J���`�+�mr�50�A9��6RN��W�kvmp��隷gsl�(&�}�������gfe�!35).cu^b��Psfה-����P8(�-8�o>:=j���*�{�Gl;�����z;u�Νx������z���z�]zb� mu9��i�d0c.+t��kw.�-�V�������=t�Y��:�ڽ���C\y痪�/�2O]��˞@=n��=�ln���g�YK��V;r��j{u��gKɟd���Ii�F�D��9���=�5�G=d��kp8��n����"���"�]\C�պ�^N�[q�SS�Hv��{nLo!w:獇�ۧ+V�=\�<�����=ixxݠ����궗u��>܏���n$�FE�5gK��6�X����b($llsǶ��ֶd���
��[�Kk�ݭ�ر����m����d��A�mp)ŷ����']��q�b�01��k{f`�=�w��">|ZjNt'0�[t蒳��2�pr�j�h�p��m����m��>�ź٬v�T�7Wl�����+��l��a�8չ{l���t�L�ju�K��u��(oG��o	�����ޞ=�]P�v�8�w�������T�tf{����}zp�V�L�%�7��ȓϭ�nx�[�h��(�oZ��e�Rks�ʗZF+*���I) �rടp��Hg�(3��Òt����B�y��d�#��!WDnv�I��6�[��1 T�d�@�^f�DK�P���*�M���`�K;;�÷;����=��m�7�u���8S>>4���R������;xB������	�*���C`��m�+N;�����xc�4]޼�p���ѻ�q��P"�ln'Ϳ�'3Q��E�O/��Wl�ȓ�Y��]R
�]���՘y �O�w�p�}Z�d�X>��Ɗ��'2KE.1���L�C���dJ�������nun�i��$�t�iCΚǣJ��|s:���х����g�1=�ϟ&"Ŀ7	d���wT����u��dM�;�h~�e�gv���%&O�`:����?R��Q��L��uE��ߓ������!Pt�1/o�jt�~SE�s˃մ���.����y� �(�Aى�\���r���q��O��D���P���N��>2�8+����6��8d����&3&�9)����w�����A����c��iՋý���
20n��;j�m6:�v�Kz����Hz�M���>[a_�ES��V{끏	�^*���[������ɖ��k*|&�'�p�4��b��τྸ��՚/�E��s�?K�\�0���p��F��{﹃'����ޙH
���3O7�r�SN2^�m�L���\�������q�:�On�p)�iGf�����f�[�[�3u�<��Ⅿ=�Q1�{ ա�x�D�zgҸ����S�� 㿣��}�%ӡ�h{�au*�@ɳv�1�
@�wy�:��؟A=�������"V��<@����Yq�D v�l��6@����oO�?*�1�m8�I�1>�Wl��0��)#7?�Qa�a�5<�(���K+�`�ۮ�ys�\�&ŗ=m���l��Tn1{l�VW��n�oYF�n]���F�Q�Vz�Г�x�oobFۀ�+.hw�(2�nvykI�î��eF��nS����~~����	|bK����M }�5Z�d�^+�_X1ި�l����^�n�Þj��)�6w��k>u�	S6��m(��7�k�����ռ���C�"K�r�H<�d���8'm^�����h�gJ�i�A� �`���� D����V�U_UT('�2!���o��������4[�M���ts�kj8�Ř���7 ����=ٵ�����4>y���I �wM*�_G�k�4��m�mk�i���ʺv��M�ɵ���$����R$su-�r�kr�}	��ǯ�j�{&8U���L���dϋ�H�=|ޘ03����S�u��|�hC��P���T�Q-m�$��H�`��1�匁�r5�#O�`7+ժ}(�r���I�Y�ƼI��.��z:�k��!��W����P���!�G��5�_x��`�[�9� ������p���]�Ӎf�@PΜ˾CC�9�S�/��l�<9��j|��4 ��pG�@���jy+�^ycb��S�țÂ��PwR��OxxʐH:��`ۡ����� uܓ��×��iܵ#E�0�Π��b��|/!��+�s��:���0�H u�� O��]��/�4!0Sp��IBE��,6�L8��r�'�*&(��=��ohf;���۵cg0z���/��"��9/F���bH��B/���*�s������W�d��L���r�gGÂC���d`4��]�F/_{[�N{&�z�܊��"d^����b�d=����2�,�����+7����4��w�T�=M�D�3"g�@�($w��D��x��Y� D⭟=�[�G���f�߾8f��䬛7���>:2f({[ �+�uf�yP�ya���[�3�h�����z(�^��`���Jh�D:��V�Z�sh���(-�т�l^F�0��J��˹��LM]:'QAP���>��Z:1� V/+�o)�&�_�'&��-���T������0�A�o:f8�sU��z�� Ly�����Q&'=6o(���B!0w<�d=��H�k���;ro�f�x�6��9N�����5s�N���nt��n��f�7X^��a�ȝ�7V�尼5�v��[=<�L6�	w�:I)
��l񺰟���*9�����><��ҰF��x��5�[��VY�.:��[�ob�n=�f�6�)o���wy�UpoJ�1��HT��x�T��B���ʛ��2[2���dS����^�X5<�k���^��<���`f�F���	ǚ���#�؞ I2��I�̙p|O�N�z;�,�襾�D"|��0S�
��`�(6��\t�a����5 }�{&�<F�ʹ�'��s-A��y�t�fx��q]�N}�H�Ț�J�;̹h�$�Pw˞q�r�5r���qvO��-P��r$�j� ���ǽ8�y�J��c�p�
;�jz��:��v{z���!߰�@��8P���j=E���M �����mv�0�Gb��7���_x��$)�_o�?q6�κ�ÐU55[j4�9�T�7��̸,�(�2I�qj��{ �$�>�"o�d.��nX��j���Y���o�B���А'�froܸ���0I5�W̓�b!���L����Ͳr�Q�݉��6
{�wg ^���n��tۅ��U�ұ��8��@e$8`v����c�â����#�o�:�V�i�7xά�̂�Pu�]��&l��&�Y�y�54���,V ����/x> o�\�����#�;���N��,�v�>p�<'&��i}l��;.�o�p�������C� �c�W�O�
*�����DS�Vj��/]���$w��S;��Y��x��ن��Q#����T¾D��M���Oh�k��B��dx�o#�V*�[���A�<����b�����Զ���|�����������>��7�jHz����ߟ��-��L\����!nRA�>�B�o�G��J�jE��N�XL����Cx9��YBi˘�Q�Ǯ�zx)+��(� h�z�m�w*�W��;?X��d����`@��BdnZY	���-�Q=&��Q�0T�W�0"�ֳ��L_��jL��̞p�Iz<R� ���-��ZP ��wt9J�`�g�R���m���oc����=mo���a-qd���l���W��B�����J��]*|�B��H�'��׵�A�a=�(�g@u�ecQo�!X쁙H�ݬ� ��#�2,����,����b�sbu���_9���IC��H�d�hX#(*�\`^5w�ٙ�~e"=�,���8+rb��������ܶO��7�)���FFT�ЯP��`��v${VW�ý���-�Q�+�9�����Wٓ;F�Fer�d�$��lܴI=V�J����هF�D�ś��q#�X-���q_P�)�1�X��<���+��25~բ*�KG�$�Qo�|6�˕���©G�^R�WmՆ���0���F�p�#�n7q�̒����{k!s�q��� ��q�q��J�;5�X�Xsa��k���pt�c�'J�O���-��&�M ���H�x��2� ͭDĤ�Ɍ֚+�fr�	�*�)p̋V�٢�X&��>��S��g� sW.q����_6{�f�ʃ���6�ҽ�]�KW<��{�]fG[SG(,�s|�U��4� P�@b���qݞ�o#lo�,G�.0��ϙ#�|����fd�*�@F���ى���s��.4���{���W8���$�FE��wK+B�J�N��}��\'	E���oeBm�*����,��k`[����HHY�j:W�ˮ�D)���O�2�!{H���s�䣺g�h�(z$�	L����#���
��'�4$q^/.,�CΌ��gɟ��������~U#g���&�i0z�P���ⷔK��#��0G��"��R�0;fN1�M��$2�g�u[Z��Ͻ��)|߷��j5C[*=TǺs�q���&т�V��x�M�շ��rC��&OxJ��m;;�V�>^�%� {i��f�(g�����$f4�ѷY��ݜÖ�7�P2%���j�T
��ڝ��e�4P�Tc�k7����}z��{O�3�6�N�-�W5XX�������	�`�
���s\9�:}|�A4�o����O����8aҔs�)%�Ւa��:�\��1���C�y�}hxA=Z\W��T��kd�@��������	���4p_�9	�POVv1�9�jՕ�:���WƘy��c����Bx�]�B��D�p��+�˗0���g)���9�'�<=�\_=�K�5`oZl^�a���)S�mi�|9��3���L�����"*���b����V�ǆ�S�9�7�"I�zP9�~��S���F�M��-d\5��W�zSht<� ��ȍ$ji�&�9&�w^'ċ���ۇ��Y�=&�?�D?N[U�wP��PTeE��~4V��][�כ���Yӗʒ�| 3 �1�z\^$W /]a�$�]lI�;�7�	%�#k�*����FNu/� B'ib�8�]��ګ��[S�Ζ�g�u�h����X�Q���h56���_����H�%w;�ۮ�=ۘ�z�.��y�t$�셷7=�Z��ݛv��x��WhKn�F�Z��Ӆ,�Cύ��n5�f��oo7�sӞ�W=��q����{�ϗ�����=��#a���(P���p�YV���%v�*�#w[��B~`C=/�Xq'(� <+TM�����x���*7�㘘C��=�A���b�_>:�:k�aa�`�:�e���^guǨ��x}�J�2]�/��skU��fP����(�������[?�s�r��. EZG-1�+\�B+���ꉱ�"L�a� �C�[��3����6��=�j_/R�d^z�_���j��P��Xׯ3-��l���Q��~ߧ�)}'�~`{W�LS�J�,{��?\+�����$pUI��k�0��k�(�������ҝI���e���ޥk�vJ��b��ǋ��M�����]FW���8��& �"�<�zsg2�Ĥ�T��T&�sk�Y���I>Gշn�?�W��1����w��n�3��;F	�̚%��	!x�שʇ��F�*�%T]��g�'������G��*˴3ػo��Rg�C&�_bk;�9���&���x��0��y)^.��N�9ص�0��D���n���޷O��������Y�% ��}�~���?�X�����$�}�{K��V+(��=>����O�o�v��-� te_Q*|��L�N�3���>�y��Q?��+��Ͽ~��N��k�`�|������)��@X/Wc}B�*i{�/��рqr<�l���.��3� U�3�Z���1_�����
C�96���m�ˆS�����P��i��N�0��o�P�
ڏm.1�&�>�֯���?e��Yg},�(,5��XWL�GooҾV%�q@/>z"�C?�;�%3[��*ϑ�G)�Y=�,����z]�bDz�p׶��>�����D�/��ϟ̛��v���ūjx�ḶZHfaZ0���Ń��Õ�b��ݽ�������'�|�nv�����K��R�7��V��O����*�����j�n�
���������WM9���GZ:�������
�}���p�=�P��m�먨����嗄�a�vR�E�DY'�����Y4�h0v.7��3��5#g��H�CH��+eK�0qX\6�����m
J'mea)4]���&��ŗJ�3��	@e�8�ة�������]�+��p=.�(�H�ZN(tZ���s��ͫ�!�'�z� ���7�f����F��] L�z��-k]���Գ)���K�t_�Ӌv��s��v�nIZ�a�.8���lx)&�VW�s��G���.a[)^I��4Ui�Kѣ��K0ޝl���/6IF7�Kg(�{�\ꀥ3�ga��a�T��KxIU8G+.=�G�������b��0��aA��$�I[h����k��I�tvN��n������oa}mƷo^\�g����h^]rc��qیW��7^�Zy�WIlk���F��\I�d��n�#X<��ѷ���t��uf�+�t jy�F��dx�4�l��ծ;	^9��F��������{=�W/Rq��b���k4q����]v��s��X�g�w�DyӢ�gu��joh6��-�u�Y5�7k��k��1�lI�k;kv���۳ӽ����y�;y��1��� g����c�d1�\�t�K�٧k�`�r<��\��[����jd㱴g:u�7+�l��m����ʨ��ڦ.�,��=������n{*{b��.�L��=q�g�y��mn����ic�&[�g!Z겖��cdM��1s��������������8Mē�0f��v��=mz�͊��\�y{)�ݺG���;�x�k)�w5[����;h\��� ��>�cu�9�5jSS����/Z��9��x1îc��!��Svv����{�z��_�|��F���T3���ʊ���t̛ݭ�z�l��	�goV��-|M�L���P#�B��_���f�!�|���ZԋS��{�Qx=�bc��[@��6ZWA�Qb�*� �H�������"���@okjL�^�B��;��P+ހ����A�$\w��mo� �8 �?#;;PARp#�SZ�m���W=��w�����i4��5�Q�e�9��&�(Z ��P3����ӝ��
�_��ܕ^�Ag��E
�9\"�%����s-�[u��/�#\hhP���P	z<Yd���4%Ggt:��I^�2 l/���L+�!"��݆UV�[R�T^�5��=!���ߌ�nĥ�2�G��<S��@��°Y�6ǐi]�t�[��؇��ƙ�՝����>~߽��e��^ca=G9{�E��˷[�P>Z�6����z-�����a1@��qu���=����,�m=�l�j����G����u�8/�w짻�|��ɗ���̃ג)^0�����"���q�׋w��p��ec�S�l�'!!.4��woQ���H�k�_�L��v~�ށnPv��{a�{��a86ߥq����w�~n��>A���ι�e�`�Xm�ɼ@|�}V�(=-G0V�'�"�8銽�h���z���ȇ�pU��e��Vn���U��"�9��]O���95�=
$���2��Jj�u��0���W����=���ŤU�)%�B2v�VV�6���k�a�����,�Q�<��F/�eC�P}dzߦ{h\x��
	�d)�D"�M��#��q�>���U����΢�˅�3XL�0���ಀP�o<�JJ�h���:�z��v��˄
���۹��,����JZ�E��{H(%1����Q]7^��ʚ��N�ё�Sa��Ttl.�U��6�{����Mk^�3k��i:�yZ��VT��(2U���M�`r��N�,�@��
J$�9��DpW�&��h5P]��;��#��\e�p�|[��g��8O)����i����x�ㇺ$P���^8�8Q����k�Q�6�d���h8`�FOx'��.7� !�5�ܝ}q�kQcI+$T&��,Vv�O]1�sW�����p�&+�ZԺ���i�|5����ɈW��������R"<p�lo�#�o;'�b3z#�����5��*4Aި�`�9{_����h�[���}V�F)�6'vj��x]������߿��w��8>�=�+G}Z#�c�y���绵2L`�U��1N^��Ĥ�<�8�Ʃ�.w�(/�aɺ2�d�n��w��!��cѳ����~����9�R���H�n����!x!�}�Ǉ���Y�J���^����a�r��n�S1"4a�Y�W�;��D��9l���5�<=[4U���3��=B��@���w>���1��Ĵ��)�Gz%���9��v�cbvb�`�U�_Yqѐ�0�P���z���x���{�o�i���lk�qC����ާ�zӶ�-H����GgZI@3���4I�DɍG�v����C���mj�\e�u�Q�np�����^�'�;���.}2��!P��*e��X���%,�x����m�Z��tk��=k̥{S[��踏��J.���'-��U���Y�`��j�Y�6���o��fH�xM{bs�?lnL�q9��S3"�5�To���Ǉ�5�*잮Hv�(ʫe��G��ٙ��|�Ġ�ETid��67�/+�QrX��E�iR�{`��JP��)�-,�f���+6�q��z��O؂��,z7s|��W��l����5�o�f�U�ܞ�i�X5�3j {|`�QЭĭ&��8�j�W�	� �G��t��ٶ"�Ъ�]�U���רۏh���2}�_L�;I��������ǺL��g**�,9�37K�䖮�.�-�y���itHY��Tl�sŧnf�ؔ�.ͩC��pr��cGK���-���
k�wd�|Ύ[�6�4h'���ln���Lm��&N���c��/`k*��;�&�h�`0!�[M$�f�{%���W]��t��"z���H����_'�or�ц\;�3�ˀ�֥���({-fh���s�^=$�Q�f缪Q��T0�yƻ��xmQ� 45�Г
&Y��͛�d�Y>��y��}~?��y7�A��o)f�A�!��Q�� �@����t����h#@v��bͪڌ��]�^pJ�����9�v���y��k���v�U=���3]�ݐL	�Dތ{�e#�8���0�VW�CUC�ح����/"�o��My-ٷ�l�g�Z(O�>�xFպ��K8���7��0v(�/���㗎����u�hyód��N�Z������46LeǮ�l4�[����s�3·W�E��g^&;��؍�6��sMwo������T�I�߳C��c��򳏘M��Skkim�մ��gx��w]gBn�<^溗-,[�Ӂ��Ƭu�. O��>j� Y+��ᆐ�����pwMB������>�s�go.o��p�W�W5]s��p��%�p�1��Fk��_�x���w{|��3E0L�}t�Wa�wK��Q����#�[��mH*�w=�`���v<�	/��#�t�w��|بzw�6�w\�;(�Qv�$8��o�����Dx��ɗԟu+�b���74��I�
jd!p����C���frN`���7����tG�u�g08jV�hGXg�'��f�X��n���ێ��iӖ,��!�c_>	�}���7�To�=��˰[�S!�� �Ka�Qd ��!�����1���g�O�+��K��z�"�`�谳��z��m���b�	�0��J��4n��ɝ}����^�l����ݜ:�]etw��XHLV{���<�o+�:�BǺ�4͂{.�͉&)�\sl}�'G[Q�����VCn.Q�}U�F�"5ꉚ�ݾ�2.v@�X�7�!0� �A��SpE��	P�N<��J��L����TՄ��q\"E�#�3&����W��]���^�]�!�~�;O=��gFx%����#��N�KS)����^��{à�d�H0��AFkݙ���YC,gNW�ȍ�q���x@�Gg�\za�3�^"��$�F:�)�dlJ��F�6�H!
�F�tUf��pk7�ݮ�F.�sŭ��Ou�C\<�\g�,a4lj���ۭj�����эg[&6����n͝�y����[��BECL�o��A�\����_,�=��ж�ce�^�%3���ն�ŷq�{��yGm�2=�61���b(���*{�Y�b�����R!s��o���j_v����~�N�%���;i-���BN���FF�#��g�끳���3����ㅍ��g��5�
�������U�q��ٞ�QȦ{#��I�6�3��º��8w��[eM؞������;���'�㕵�Ws�[�{�^�e5p>j�p?���/E�b�ƨG�u�z/G��d�o��u�*����Y���5�eece��s"Fi���T���ݳ��Ǆo!Cp\� ^�k��:����?��tno��f�;����s4a)�k�j�u�Xc�����z��n�����΂�F{H�G��=.ze��_i�J�:��*�Þ�sMXs)]�����ޒ�n���n_6ؿG(Ge�Lj�n��W�|���=Yp{�/�}��A,���B;�w!��$q8�!( Cl�R��5��QsG��M��=��?���
�������h����l�2���K�W�BK�}s��i�	�F�;
E�"�o�:���ΓS��g������(��㾣[RM�G?v{�7k��z��`�M|����hb��|FL�-f���Ie��(� ��;�3�b&a��>s����)�3�����
"�?f5%Bm�ReV�zj��ͤ��j�=�n�\�NaC�5����*w�|A��6Oy���]+*֜�r�w�3�~������yoGY_eR���ɇ���9<�hgP�:2z[��b�D\�u��S,�^���Þ�;��{���_`�9�~�6G��{�����Erbk��,hߗ����5��6�<sԡ�Pg�;���s��[=�E�o<���#��,pa���O�u�v�w���:y��v�و*'Eg��S���Vܼ�e�@U���͉s�~'��G�"��o_Ev㚐���쎏CdB�O[�}��:�yX�]���h��Bj�*(���@P=�Vw�:j��> ����\~z
;��?#���a��a��E,������ ��8��������?7}�s��8:|u̧4`��6�4�G��ڱ�3��wUϕ!�fgfW?��
0�*�'��N�n�S��Z9��x����EI���f�h�ݰc�d��nd\�'�+��=��٢"�p��#������F�%Z73,����-3�V@l	ؿ�u�XR.�w��
w.p/���vȋuxD���'5Ӟ)�RU=���SէT�T~��#,^������,���
zD�	�VK���듾=��op�]�����E�RU^�2㿶��9r�=��Ժ�Mwٕ��%p�Yao>��箊~�Q�X�bR)���G��g2���0�s3-����e�zX�G�D����wh]�z>��?���=���gm�]�v{=�`�p�1
Tz�]� fl`��w]fx�a�=��~���$v�'���؎����ݛ$�W�#�Д���yyU{��ca+���Vހ���u�8w��"��I�O�l�t���.+)�')�����}���\� ���^˳�Z)m�_H$��+{vcB�X2�ћ\|` g<�y��G1���p,希P�E��\_����,��<���Q�0�z�0��>���b����f�eWu��J;���B�eE��@\�B�q+��u$��x7W�5���U!��~�zki��a�F�c���{u�=�:3����q�֬�MV���23�c��vQ�� |��!ࡕ�z�\(����n� r}|{��U�̙�T�S{���h���{��.к��&*'�oA{�L�S�Ǯ�Q&r;��r�d�7�bP�zm�懡p��`J���TY\+NSor� ��V�pM�͎݊s�iT�-�SV7��B�lq\��/�Vֱ��������$��,�ه)D�����Ýi�N��(:� ��;��2���O��-E��y�.���X���p�P�mCY�4����71K�ҷ�K�su�V��v.�b���6��55�i�D�KBVm���ڵ��F�Y]#���l�z�yg��u8M����`�/n�rciq�9�9�t���e�[y������a�v�q�����̝��n�Q��fy��n
�1�,�Ưg���W��e�۞���S���gq�{=���OU�6�̉�a��u�ٷ62���`��I��n�@��w��g� M�.��2�nAZ�)��	���v�하+n��+���ίX�z�[�g�H���]Cس��:}v�:I+�g�N�s�l<��F�6�._n�A���z-��:�E�ہ�ՓN.�Y99����ӻ[k��B���_]��q�Fꍇf5ƺW<3r����p����>�97�m�N�o%�۬.:<]��=���}l��)]���OL`�:6l=soQ�j5|��O����w��?����V�3aí����;��չR��p'k<Q��8/0j�q��;%���8��K��3�h���c'j�V����q�ӛ���vzmٽ�;lOmۨČ��hsl������~~����ݻZ��=��DO���a�]r�{@n�����v�6�b�ն
��i�0�٘Y��1�5���%FO�� v�3#��׬>��<,�tn߯��m����k��BnUZZf��o��oܶ�������d�T���mK�Q`����$�������6}{�Ì��������y��˓�yHB�
ʻ5�Q|̇G�#�]˩�a�n&".��>��{�6��[ﳑ)��]�V�5G&<�a�!�n��4����ݝ{��m�D�\MpɊ���I/9�.D�H�M�#t�����`ov؊E_�RP �!6�)C�7;�5��zi������N�������E�O��!>�i"sވ�ߨ��x< ��K��K$��3����s�b��ݏd9���O�*MT�0"f��ii8�dx�'��ff�dT�d+�(����Qǳ9�������t��.�hm�i��.�3^3�$c�g\c��Y/�7���}�?��Ë��/��Ga�8��jfO��;3*�}������w���T��^��63M1՞8W�M����z�=>ڌnߑ8�Uݹ
�77Q�)w*��n�&g�&`�p�t=��_��������t�7S1ʠ��o������\,�4vl�z�mw�򃺎��	��ӣq���@����[���������7v�h����A)"�$&� �0�6X���g(���� �<�H��q���C��8�FǗ���j﫯�%�>�Gd�Y�W�;���t��ec�Ce�Hy~��ڮ'�n�����vbi$����e*ћSCض6:���`1�ojMP4٪_jJe�B�!De,�FoQq���ڭ���x��������j{v�N����]J�9�e	�޻n�fzgs{s[km��#vK��Ǫ�u�v'm�P�3v�g�غ�����qIb������j�߿v��mF·��y��������f�AH�<3r�d�ZkpהI�"��f�NUd)�FӇ��Pc��V9�s9�\y���P���f�4�+�B���2��&D'v�J�|'�dc��&��#j�ܞ��Y��ǧ'�}]���f�����_8E�4�0X��p�e�Y��gq:A���z�O�q��c���v:��	�wv�d���ϰ���d�'/W6�
����@��kލ��^5���Cn�E4Y
�/�;S���S�b������ϔ,���]g�ǔ�y��Ps#nz�����=������PN+h��y��=��a��ܗ��|���}폳���L��� �
7 =�FOvL�>&4q
9
s�ÅװF��	�f'�T��[��O��쑩ߒ�q�9�=>�5�m��T�v<̖at�9�q�e�9��Q�����z`wu��S��.#�g;��1q�Cƣ��e��i�u�S�����_T����#�
����G���m${��T�B
6����=��A=}��y�_��(���^�Ics�Wc����w�V�ׯ�=���܄_ս�% ��O͟����Ʉbi,�Np�89w�6���t�/T_;�>�U��-b\�ZEU=��C���H3z���m����cy��紮��Or��=����&��{j�N S}���b��J�%�.Ȧ�fp���z1�%��������V�����B�V�ￂ���w٘�?t�*~�^Ѱ�n���q���ttS�Açݱ�9壩���Ud".W�_g;
}Y�C��c٦AB6�ϧ^]S���Mx�[z����d#����y��\b��Q��ȗ.�]ƽ����V`w��n�]�,�&�K�^(���}t�:7t�B���l)�H0cqsrokj�vQ�x��ù�u��fn�ϗ!���Vw]�6l<7�q�jm@̜��!�;z��6��{q��i�PP�!큞��:=Q��@�=ӯ�Dm�fBm�����ˣ�q�H9�����͕Z���_�,����<�w�Å��;���Wki��07r�צPӞ~͏�q��(w��r�G�\��=����b=!w gs���ѿx6���Z��/[6�`8n�����Hoz��P�C��TS�Q���Zs��mV��Z��Hԩ��L�]v�5f�f�q��f��'����c׫�yF᪀��J�Բ�s{����yz9�z���]���U�l�9�a�2����klw!���p`?FP<;J��r}�_����C$.a�[hv��S2�n�A��=7ck��� �����gr7=�]0���3:���뷃�QN=w���[u-'Ͻ��:����(�[���\?�+�~:��|��ޙ��F�C-���5VCn��tj+�r�=�6��͔���3�~c�MV�\{q��ڇB@'pԒN=�7���/3.���4�+7V ņ�8��1=��1���ʛ��*Rgeb�ރV�ؕۋi$S
1w}�$[|� I�W���o4�t���b�ݘ�RK�ب���tI�N[��WLMc��.����kf�z��4���7�yNn%]a�z_���x�%��]�iv���9�;N	�)�:���m�ݵ�q2�U�:�K9*$Wv�X�,K�XW�8R�Pj�#���@Y�[ގ-T6��-�X�%+��������X#=W��]��KgD��J���>��;�zxh�sO�敋��g��y����(�!�� ?���i��L>��Ѱ��>����U��D��<����/;����q��x\�E�RQ�b}�ev�F���Y�f0�\' vwl4x��8e�֍�7����|����%��{J�� U%�2y�[q<�������U�z"����7GZ���!�ӱʶ0���0fgu�n8��
� jG_O.U���r�wfW�t�O${�,Ƙ]N(L_�T��П�
�u͂�!������R�혯wR�]����AOv�/�� ���wVwe-�TH�pM��N��ـ��*^�h��*z�pޚ^�f��'��+�l7I��%���_����ӛ�w̍���Hy�q� >]Θ0.Ž�8&a1Xy�z�i"O�o]�=,��ܶ ���^.nu#ԧ5ɴ�:�d�&;7>��A�Z�S�WJ][��"NǮǸf
"0|�vci����V��������;���5>鑐��͂���������#���nO,����\�h�d�"�c��?o����䧝�~�Su����)1�Zd�h�5X�8���������|��\c��r+v�8~j��)��f5�f��/���qo�~��i��է���Č���Mx���&�O���75�醰�Ϊ!^��5��pf*=}?y{r�����io�w^�nߞt�Eq/�7�:�j��K��x|3��a������� �I
�ۨ��1`�$v����j�7�&��ѵ�\�S��?~y���>G<��Y����2���^�r�UV��ޫ�鉆��ۇ��=7C!��G7��8�';�oq ���{�$u_��i2��u��u���s4��jCίڿ2�v��ً���n<KU����Z4���ZQ)/!u[~<yc�VY�F��]�8p�%H��*`����y�H����n�d�?X�$-0�&��x��b�Sr�g$�({��zN�\��p�Ob��ͥ�}�QU`X"3���z2��p������vR�`�}��퉂8o}e��0��<��g�O)+3��ǐ���2�o|�V��f)p�Q^�C���d��Cb.�ڿ�1c���}��z���s���\�ws��Ꝁ���^�!J��V�̈j�[	��z8�g`�W�Xf^�
�T�8Ho�uϪ�T���n_x��-�n��{6���gcI��@G�P�qrP{�����_hM6�J��2�X��~�>���ܨf@#����79v��Z�qf7��j'B�4�$���6�,��5�����������7���ō��\�[�-�&�:�����v��v�Fƻ��Q]���8�	�ᛇLdm�g��;�qB4U)b+�Y�A��ݤ���7;�F�2��)׋%�)>��P�����3���X:h@�����o�c**����[����mV[��ȸ��Ո_\.�+��R��e�g�۾;)������I����2�Fyq� u�)ei�Jp�	��}��-��9����=�v�O��z3��ez��0��S��Wv��Y�]3�u��Yu������V?m�-���:h�.���k�`��]~/''��ί�lB��yP�l�j!�<��7}�n�|�S$��xпD��Q|�S�p�noMML��-�������&2{��oM-ݓT��$����uL�l�[�($⸋��q��wؑ!��
=Z�����/ ��~}w�}s��[�^��4�αQ0���h�;��ǽ�Fm�eWe����l�)���о6F���=��O����:aI�� �I;�+�>�x�ѭ�9i�}�þY^k��.�������3/���
�����Y�^ E��� ~�-/C���l_�qv�w�����G��2M�$�0� CA�)�m�q�"-��n�V���p7�㦅ˌ�A�wGt�`w�1o�P��ݕ��f_
(�g�w�z��t&/˺��``�������\�o�p�ʽ�c���Զ�����tk{7�~�<��X��U�����7@n=;�;etZ�R��������K�%��m��m��S�-��O����ٳսf�i���ZQl�f#w��ٍ���]I����j�)g��3vG!A����5ZŢ�ÖZ'�ȋ��=�~28���ǳ�;��;�	0'4�O{%i����j�֫��ڮe�V���JtB�����h��UTY�#,!	$�	O�>�I�y����0g��t;��\,�w�f[�N/"dr��a�d&�Q�!FbBBp�
 �$ ���aHI� I')è � $�	��@�f"���P	$a A� HH�$����}����1;�� r��\��=g�H�H1X�w	��[b��V�k���-�v�O�{�ͼ*�i�ST�Q��0�z���<���ok����&��M/crί���i�]��t?���c^�nzU�Sq��T�u���칉�c{w���zLgF�����{\b"I#Ȝ����<x��+�4�����$���;�}0$$��#$!$��B�J����Jkn�j�Rrj����(�.s�*<:LG��/��1�}�nɧ:�ؑ�됉$�>�{�'�Sع�X�t?a�0��i�i�2l�0�&��!C��&�Է��!F	=�:b~o��Y�a��͋#��\�Ȧ\~CΞ��|-�OzzY`{?������&���@�A�!b	&�	$	(BN�L>sd��L��XB$�(��!$��	$ � 	!�a!��"A H�ی��d��$���z�.f�W^/�6���Õ�rO�B$�9$Ɗ�qb�dUk�>�s9�5:�������%̗'W�S�2�����r��XŴfEpԘ���k�³9�o���8͋�"I"��u'b�o�;0�Oɫ���Y��f��sx���#;ƷX�d�av!�鳾�_R�̣�S^c�b;�JpM�X�Z�.��ͯ��O+�!IM�V �#��;�/��G�
Ga/����ǘ�q�C�~O �v�e%
20�g��		$�ú@��C�>��}��<I��ì=�J��Ə�~�i�$��lp22�>Tā�؇�va�$$���<�pn[RФ�b�O4�C�ǬHI HBI@@C(}�C���@�rIۨ��(&��?m�����~%�>�����w����q/�+��p��i��GH|����w3�d�iI|���a��{�I$<�+:���C�����_�eI>w�~ux���\Z���6�z�T�����JxEg���{'�4�|C�C�����U<�BnT���^UM�bg�y��@��Ci�p��&�%��	O�D�dI$('��0�;���SkF�n�	�N�lS|����Vɢ{zI���' !O�����p��QB�.0eEL%x\L�Z,ka�UFJ�.��>i��I��M�<��)OO'} �3a��L�y���ϴ� BI!JO�w�xE)�\�`rE��~�G�02|���6�4r68���t�f����38�^潽��!��:HC�;���C�<��!$�����%��0<�!c�0jM�!ԥ��`��:B�H|����y@�q0L�{��{�ﬖ&s�>Fm��G����e�S�o7���)��~��i��$�����ܑN$"�� 